`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:02:53 02/25/2013 
// Design Name: 
// Module Name:    fowarding_unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fowarding_unit(
	 input clock,
	 input rs,
	 input rt,
	 input wb_ex,
	 input wb_mem,
	 input ex_out,
	 input mem_out,
	 output sel_0,
	 output sel_1	 
    );


endmodule
