module uart_tx
  #(
    parameter DBIT = 8,        // número de bits de datos
              SB_TICK = 16   // número de ticks para bits de stop
  )
  (
    input wire clk,
    input wire tx_start, s_tick,
    input wire [7:0] data_in,
    output reg tx_done_tick,
    output wire tx
  );
  
  //Declaración de estados simbólicos
  localparam [1:0]
      idle  = 2'b00,
      start = 2'b01,
      data  = 2'b10,
      stop  = 2'b11;
      
  //Declaracion de señales
  reg [1:0] state_reg, state_next;
  reg [3:0] s_reg, s_next; //Numero de sampling ticks para hacer el oversampling
  reg [2:0] n_reg, n_next; //Numero de bits de datos recibidos en el estado data.
  reg [7:0] b_reg, b_next;
  reg tx_reg, tx_next;     //Buffer de un bit para filtrar posibles fallos
  reg [4:0] auxs;
  reg [3:0] auxn;
  
  //Cuerpo
  //Registros de datos y Estado de la FSMD
  always @(posedge clk)
    begin
      state_reg <= state_next;
      s_reg <= s_next;
      n_reg <= n_next;
      b_reg <= b_next;
      tx_reg <= tx_next;
    end
      
  // FSMD next-state logic y unidades funcionales
  always @*
  begin
    state_next = state_reg;
    tx_done_tick = 1'b0;
    s_next = s_reg;
    n_next = n_reg;
    b_next = b_reg;
    tx_next = tx_reg;
    
    case (state_reg)
      idle:
      begin
        tx_next = 1'b1;
        if(tx_start)
        begin
          state_next = start;
          s_next = 0;
          b_next = data_in;
        end
      end
      
      start:
      begin
        tx_next = 1'b0;
        if(s_tick)
          if(s_reg == 15)
          begin
            state_next = data;
            s_next = 0;
            n_next = 0;
          end
          
          else
			 begin
            auxs = s_reg +1;
				s_next = auxs[3:0];
			 end
      end
      
      data:
      begin
        tx_next = b_reg[0];
        if(s_tick)
          if(s_reg == 15)
          begin
            s_next = 0;
            b_next = b_reg >> 1;
            if(n_reg == (DBIT - 1))
              state_next = stop;
            else
            begin
					auxn = n_reg + 1;
					n_next = auxn[2:0];
				end
          end
          
          else
			 begin
            auxs = s_reg +1;
				s_next = auxs[3:0];
			 end
      end     
            
      stop:
      begin
        tx_next = 1'b1;
        if(s_tick)
          if(s_reg == (SB_TICK - 1))
          begin
            state_next = idle;
            tx_done_tick = 1'b1;
          end
          
          else
			 begin
            auxs = s_reg +1;
				s_next = auxs[3:0];
			 end
      end
      
    endcase
  end
  
  //Salida
  assign tx = tx_reg;
  
endmodule
