`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:38:51 11/14/2012 
// Design Name: 
// Module Name:    program_memory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
// En vez de hacer una memoria de 8bits y tener que avanzar el pc de a 4 hago una memoria de 32 y avanzo de a 1
//	entonces no necesito el sumador +4.
//////////////////////////////////////////////////////////////////////////////////
module inst_mem(
    input [10:0] addr,
	 input clock,
    output [31:0] inst
	 //input salida del hazard detection unit
    );
	
	integer i;
	reg [31:0] memoria [0:2047];
	reg [31:0] aux = 0;
	
	initial
	begin
		for (i = 0; i < 2048; i=i+1)
			memoria[i] = 32'b00000000_00000000_00000000_00000000;
		
		memoria[0] = 32'b000000_00001_00011_00010_00000_100010; 	//SUB r2,  r1, r3   -> r2 = -5
		memoria[1] = 32'b000000_00010_00101_01100_00000_100100;  //AND r12, r2, r5   -> r12 = -5
		memoria[2] = 32'b000000_00110_00010_01101_00000_100101;	//OR 	r13, r6, r2   -> r13 = -1
		memoria[3] = 32'b000000_00010_00010_01110_00000_100000;	//ADD r14, r2, r2   -> r14 = -10
		memoria[4] = 32'b101011_00010_01111_00000_00001_100100;	//SW r15, 100(r2)   -> r15 have 5
		memoria[5] = 32'b000100_00010_01100_00000_00000_001001;	//BEQ r2, r12, 9	  -> Pc = 15
		memoria[6] = 32'b000000_00010_00101_01100_00000_100100;  //AND r12, r2, r5   -> STALLED INST
		memoria[7] = 32'b000000_00110_00010_01101_00000_100101;	//OR 	r13, r6, r2   -> STALLED INST
		memoria[15] = 32'b000000_00001_00011_00010_00000_100110; //XOR r2, r1, r3    -> r2 = 5
		memoria[16] = 32'b000000_00011_00010_00001_00000_100111; //NOR r1, r2, r3    -> r1 = -16
		memoria[17] = 32'b100011_01100_01000_00000_00001_100100; //LW r8, 100(r12)   -> r8 = 5

		//This instruction is used to have a value to load.
		memoria[18] = 32'b101011_01100_10000_00000_00001_100100;	//SW r16, 100(r12)  -> r16 have -1431655766 TAKE CARE OF THIS INSTRUCTION
		memoria[19] = 32'b000101_00001_00011_00000_00000_001001;	//BNE r1, r3, 9
		memoria[20] = 32'b000000_00010_00101_01100_00000_100100;  //AND r12, r2, r5   -> STALLED INST
		memoria[21] = 32'b000000_00110_00010_01101_00000_100101;	//OR 	r13, r6, r2   -> STALLED INST
		memoria[29] = 32'b000000_00000_00010_00100_00011_000000; //SLL r4, r2, 3     -> r4 = 40
		memoria[30]= 32'b000000_00000_00110_00111_00001_000010;  //SRL r7, r6, 1     -> r7 = 6
		memoria[31]= 32'b000000_00000_00101_01000_00001_000011;  //SRA r8, r5, 1     -> r8 = -3
		memoria[32]= 32'b000000_01111_01110_01001_00000_000110;  //SRLV r9, r14, r15 -> r9 = 134217727
		memoria[33]= 32'b000000_01111_01110_01010_00000_000111;  //SRAV r10, r14, r15-> r10 = -1
		memoria[34]= 32'b000000_01111_00010_00111_00000_000100;  //SLLV r7, r2, r15  -> r7 = 160
		memoria[35]= 32'b000000_00010_00111_01000_00000_100000;  //ADDU r8, r7, r2   -> r8 = 165
		memoria[36] = 32'b000010_00000_00000_00000_00000_101110;	//J 46				  -> Pc = 46
		memoria[37] = 32'b000000_00010_00101_01100_00000_100100;  //AND r12, r2, r5   -> STALLED INST
		memoria[38] = 32'b000000_00110_00010_01101_00000_100101;	//OR 	r13, r6, r2   -> STALLED INST
		memoria[46]= 32'b000000_01000_00111_01001_00000_100011;  //SUBU r9, r8, r7   -> r9 = 5
		memoria[47]= 32'b000000_00010_00011_00100_00000_101010;  //SLT r4, r2, r3    -> r4 = 1
		memoria[48]= 32'b000000_00011_00010_00100_00000_101010;  //SLT r4, r3, r2    -> r4 = 0
		memoria[49]= 32'b100000_01100_01000_00000_00001_100100;  //LB r8, 100(r12)   -> r8 = -86
		memoria[50]= 32'b100001_01100_01001_00000_00001_100100;  //LH r9, 100(r12)   -> r9 = -21846
		memoria[51]= 32'b000011_00000_00000_00000_00000_111101;	//JAL 61				  -> Pc = 61 _ r31 = 52 
		memoria[52] = 32'b000000_00010_00101_01100_00000_100100;  //AND r12, r2, r5   -> STALLED INST
		memoria[53] = 32'b000000_00110_00010_01101_00000_100101;	//OR 	r13, r6, r2   -> STALLED INST		
		memoria[61]= 32'b100111_01100_01010_00000_00001_100100;  //LWU r10, 100(r12) -> r10 = -1431655766
		memoria[62]= 32'b100100_01100_01011_00000_00001_100100;  //LBU r11, 100(r12) -> r11 = 170
		memoria[63]= 32'b100101_01100_01101_00000_00001_100100;  //LHU r13, 100(r12) -> r13 = 43690
		memoria[64]= 32'b101000_01100_01010_00000_00001_100100;  //SB r10, 100(r12)  -> 170 should be stored.
		memoria[65]= 32'b101001_01000_01010_00000_00001_100100;  //SH r10, 100(r8)   -> 43690 should be stored.
		memoria[66]= 32'b100011_01100_01001_00000_00001_100100;  //LW r9, 100(r12)   -> r9 = 170
		memoria[67]= 32'b100011_01000_01010_00000_00001_100100;  //LW r10, 100(r8)   -> r10 = 43690
		memoria[68]= 32'b000000_00111_00000_00000_00000_001000;	//JR r7				  -> Pc = 160
		memoria[69] = 32'b000000_00010_00101_01100_00000_100100;  //AND r12, r2, r5   -> STALLED INST
		memoria[70] = 32'b000000_00110_00010_01101_00000_100101;	//OR 	r13, r6, r2   -> STALLED INST		
		memoria[160]= 32'b001000_00111_01011_00000_00000_001000;  //ADDI r11, r7 + 8  -> r11 = 168
		memoria[161]= 32'b001000_00111_01100_00000_00000_001000;  //ADDIU r12, r7 + 8 -> r12 = 168
		memoria[162]= 32'b001100_01011_01101_10000_00011_110000;  //ANDI r13, r11&33008 -> r13 = 160
		memoria[163]= 32'b001101_01011_01110_10000_00011_110000;  //ORI r14, r11|33008 -> r14 = 33016
		memoria[164]= 32'b001110_01011_01111_10000_00011_110000;  //XORI r15, r11^33008 -> r15 = 32856
		memoria[165]= 32'b000000_01001_00000_10101_00000_001001;	//JALR r21, r9		  -> Pc = 170
		memoria[166] = 32'b000000_00010_00101_01100_00000_100100;  //AND r12, r2, r5   -> STALLED INST
		memoria[167] = 32'b000000_00110_00010_01101_00000_100101;	//OR 	r13, r6, r2   -> STALLED INST		
		memoria[170]= 32'b001111_00000_10000_00000_00000_000101;  //LUI r16, 5        -> r16 = 327680
		memoria[171]= 32'b001010_01000_01011_11111_11111_111011;  //SLTI r11, r8, -5  -> r11 = 1;
		memoria[172]= 32'b001010_01001_01100_11111_11111_111011;  //SLTI r12, r9, -5  -> r12 = 0;
		memoria[173]= 32'b001011_01000_01101_00000_00000_000101;  //SLTIU r13, r8, 5  -> r13 = 0;
		memoria[174]= 32'b001011_00100_01110_00000_00000_000101;  //SLTIU r14, r4, 5  -> r14 = 1;
	end
	
	always@(posedge clock)
	begin
		aux = memoria[addr];
	end
	
	assign inst = aux;
endmodule
