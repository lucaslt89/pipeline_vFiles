`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:00:50 02/25/2013 
// Design Name: 
// Module Name:    ex_mem_reg 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ex_mem_reg(
    input wb_entrada,
    input m_entrada,
	 output wb_salida,
	 input clock,
    input [32:0] resultado,
    input [32:0] dato_1,
    input [32:0] dato_2,
    output [32:0] salida
    );


	
endmodule
